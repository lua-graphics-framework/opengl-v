module main
import versions

fn main() {
	versions.gl_viewport(10, 10, 100, 100)
}
