module versions

pub fn gl_viewport(x int, y int, width int, height int) {
	C.glad_glViewport(C.GLint(x), C.GLint(y), C.GLsizei(width), C.GLsizei(height))
}
